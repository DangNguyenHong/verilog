`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:29:51 09/20/2023 
// Design Name: 
// Module Name:    MUX41 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MUX41(
input wire [7:0]e,
input wire [7:0]f,
input wire [7:0]g,
input wire [7:0]h,
input wire [1:0]mode,
output reg [7:0]led
    );



endmodule
